module TMatrixMultiplication

MatrixMultiplication bluePill();
endmodule
